package shared_package;
	int correct_count = 0;
	int error_count = 0;

	logic test_finished;
	
endpackage : shared_package